module mux8x1_32_bit(
  input [2:0] sel,
  input [31:0] in0,
  input [31:0] in1,
  input [31:0] in2,
  input [31:0] in3,
  input [31:0] in4,
  input [31:0] in5,
  input [31:0] in6,
  input [31:0] in7,
  output [31:0] Result
);


  wire [2:0] sel_not;

  wire [7:0] and0;
  wire [7:0] and1;
  wire [7:0] and2;
  wire [7:0] and3;
  wire [7:0] and4;
  wire [7:0] and5;
  wire [7:0] and6;
  wire [7:0] and7;
  wire [7:0] and8;
  wire [7:0] and9;
  wire [7:0] and10;
  wire [7:0] and11;
  wire [7:0] and12;
  wire [7:0] and13;
  wire [7:0] and14;
  wire [7:0] and15;
  wire [7:0] and16;
  wire [7:0] and17;
  wire [7:0] and18;
  wire [7:0] and19;
  wire [7:0] and20;
  wire [7:0] and21;
  wire [7:0] and22;
  wire [7:0] and23;
  wire [7:0] and24;
  wire [7:0] and25;
  wire [7:0] and26;
  wire [7:0] and27;
  wire [7:0] and28;
  wire [7:0] and29;
  wire [7:0] and30;
  wire [7:0] and31;


  not not0(sel_not[0],sel[0]);
  not not1(sel_not[1],sel[1]);
  not not2(sel_not[2],sel[2]);
  

  and i00(and0[0], sel_not[0], sel_not[1], sel_not[2], in0[0]);
  and i01(and0[1], sel[0], sel_not[1], sel_not[2], in1[0]);
  and i02(and0[2], sel_not[0], sel[1], sel_not[2], in2[0]);
  and i03(and0[3], sel[0], sel[1], sel_not[2], in3[0]);
  and i04(and0[4], sel_not[0], sel_not[1], sel[2], in4[0]);
  and i05(and0[5], sel[0], sel_not[1], sel[2], in5[0]);
  and i06(and0[6], sel_not[0], sel[1], sel[2], in6[0]);
  and i07(and0[7], sel[0], sel[1], sel[2], in7[0]);

  or or0(Result[0], and0[0], and0[1], and0[2], and0[3], and0[4], and0[5],and0[6],and0[7]);


  and i10(and1[0], sel_not[0], sel_not[1], sel_not[2], in0[1]);
  and i11(and1[1], sel[0], sel_not[1], sel_not[2], in1[1]); 
  and i12(and1[2], sel_not[0], sel[1], sel_not[2], in2[1] );
  and i13(and1[3], sel[0], sel[1], sel_not[2] , in3[1]);
  and i14(and1[4], sel_not[0], sel_not[1], sel[2], in4[1]);
  and i15(and1[5], sel[0], sel_not[1], sel[2], in5[1]);
  and i16(and1[6], sel_not[0], sel[1], sel[2], in6[1]);
  and i17(and1[7], sel[0], sel[1], sel[2], in7[1]);

  or or1(Result[1], and1[0], and1[1], and1[2], and1[3], and1[4], and1[5],and1[6],and1[7]);

  and i20(and2[0], sel_not[0], sel_not[1], sel_not[2], in0[2]);
  and i21(and2[1], sel[0], sel_not[1], sel_not[2], in1[2]); 
  and i22(and2[2], sel_not[0], sel[1], sel_not[2], in2[2] );
  and i23(and2[3], sel[0], sel[1], sel_not[2] , in3[2]);
  and i24(and2[4], sel_not[0], sel_not[1], sel[2], in4[2]);
  and i25(and2[5], sel[0], sel_not[1], sel[2], in5[2]);
  and i26(and2[6], sel_not[0], sel[1], sel[2], in6[2]);
  and i27(and2[7], sel[0], sel[1], sel[2], in7[2]);

  or or2(Result[2], and2[0], and2[1], and2[2], and2[3], and2[4], and2[5],and2[6],and2[7]);

  and i30(and3[0], sel_not[0], sel_not[1], sel_not[2], in0[3]);
  and i31(and3[1], sel[0], sel_not[1], sel_not[2], in1[3]);
  and i32(and3[2], sel_not[0], sel[1], sel_not[2], in2[3]);
  and i33(and3[3], sel[0], sel[1], sel_not[2], in3[3]);
  and i34(and3[4], sel_not[0], sel_not[1], sel[2], in4[3]);
  and i35(and3[5], sel[0], sel_not[1], sel[2], in5[3]);
  and i36(and3[6], sel_not[0], sel[1], sel[2], in6[3]);
  and i37(and3[7], sel[0], sel[1], sel[2], in7[3]);

  or or3(Result[3], and3[0], and3[1], and3[2], and3[3], and3[4], and3[5], and3[6], and3[7]);

  and and40(and4[0], sel_not[0], sel_not[1], sel_not[2], in0[4]);
  and and41(and4[1], sel[0], sel_not[1], sel_not[2], in1[4]);
  and and42(and4[2], sel_not[0], sel[1], sel_not[2], in2[4]);
  and and43(and4[3], sel[0], sel[1], sel_not[2], in3[4]);
  and and44(and4[4], sel_not[0], sel_not[1], sel[2], in4[4]);
  and and45(and4[5], sel[0], sel_not[1], sel[2], in5[4]);
  and and46(and4[6], sel_not[0], sel[1], sel[2], in6[4]);
  and and47(and4[7], sel[0], sel[1], sel[2], in7[4]);

  or or4(Result[4], and4[0], and4[1], and4[2], and4[3], and4[4], and4[5], and4[6], and4[7]);

  
  and i50(and5[0], sel_not[0], sel_not[1], sel_not[2], in0[5]);
  and i51(and5[1], sel[0], sel_not[1], sel_not[2], in1[5]);
  and i52(and5[2], sel_not[0], sel[1], sel_not[2], in2[5]);
  and i53(and5[3], sel[0], sel[1], sel_not[2], in3[5]);
  and i54(and5[4], sel_not[0], sel_not[1], sel[2], in4[5]);
  and i55(and5[5], sel[0], sel_not[1], sel[2], in5[5]);
  and i56(and5[6], sel_not[0], sel[1], sel[2], in6[5]);
  and i57(and5[7], sel[0], sel[1], sel[2], in7[5]);

  or or5(Result[5], and5[0], and5[1], and5[2], and5[3], and5[4], and5[5], and5[6], and5[7]);

  and i60(and6[0], sel_not[0], sel_not[1], sel_not[2], in0[6]);
  and i61(and6[1], sel[0], sel_not[1], sel_not[2], in1[6]);
  and i62(and6[2], sel_not[0], sel[1], sel_not[2], in2[6]);
  and i63(and6[3], sel[0], sel[1], sel_not[2], in3[6]);
  and i64(and6[4], sel_not[0], sel_not[1], sel[2], in4[6]);
  and i65(and6[5], sel[0], sel_not[1], sel[2], in5[6]);
  and i66(and6[6], sel_not[0], sel[1], sel[2], in6[6]);
  and i67(and6[7], sel[0], sel[1], sel[2], in7[6]);

  or or6(Result[6], and6[0], and6[1], and6[2], and6[3], and6[4], and6[5], and6[6], and6[7]);
  
  and i70(and7[0], sel_not[0], sel_not[1], sel_not[2], in0[7]);
  and i71(and7[1], sel[0], sel_not[1], sel_not[2], in1[7]);
  and i72(and7[2], sel_not[0], sel[1], sel_not[2], in2[7]);
  and i73(and7[3], sel[0], sel[1], sel_not[2], in3[7]);
  and i74(and7[4], sel_not[0], sel_not[1], sel[2], in4[7]);
  and i75(and7[5], sel[0], sel_not[1], sel[2], in5[7]);
  and i76(and7[6], sel_not[0], sel[1], sel[2], in6[7]);
  and i77(and7[7], sel[0], sel[1], sel[2], in7[7]);

  or or7(Result[7], and7[0], and7[1], and7[2], and7[3], and7[4], and7[5], and7[6], and7[7]);

  and i80(and8[0], sel_not[0], sel_not[1], sel_not[2], in0[8]);
  and i81(and8[1], sel[0], sel_not[1], sel_not[2], in1[8]);
  and i82(and8[2], sel_not[0], sel[1], sel_not[2], in2[8]);
  and i83(and8[3], sel[0], sel[1], sel_not[2], in3[8]);
  and i84(and8[4], sel_not[0], sel_not[1], sel[2], in4[8]);
  and i85(and8[5], sel[0], sel_not[1], sel[2], in5[8]);
  and i86(and8[6], sel_not[0], sel[1], sel[2], in6[8]);
  and i87(and8[7], sel[0], sel[1], sel[2], in7[8]);

  or or8(Result[8], and8[0], and8[1], and8[2], and8[3], and8[4], and8[5], and8[6], and8[7]);

  and i90(and9[0], sel_not[0], sel_not[1], sel_not[2], in0[9]);
  and i91(and9[1], sel[0], sel_not[1], sel_not[2], in1[9]);
  and i92(and9[2], sel_not[0], sel[1], sel_not[2], in2[9]);
  and i93(and9[3], sel[0], sel[1], sel_not[2], in3[9]);
  and i94(and9[4], sel_not[0], sel_not[1], sel[2], in4[9]);
  and i95(and9[5], sel[0], sel_not[1], sel[2], in5[9]);
  and i96(and9[6], sel_not[0], sel[1], sel[2], in6[9]);
  and i97(and9[7], sel[0], sel[1], sel[2], in7[9]);

  or or9(Result[9], and9[0], and9[1], and9[2], and9[3], and9[4], and9[5], and9[6], and9[7]);

  and i100(and10[0], sel_not[0], sel_not[1], sel_not[2], in0[10]);
  and i101(and10[1], sel[0], sel_not[1], sel_not[2], in1[10]);
  and i102(and10[2], sel_not[0], sel[1], sel_not[2], in2[10]);
  and i103(and10[3], sel[0], sel[1], sel_not[2], in3[10]);
  and i104(and10[4], sel_not[0], sel_not[1], sel[2], in4[10]);
  and i105(and10[5], sel[0], sel_not[1], sel[2], in5[10]);
  and i106(and10[6], sel_not[0], sel[1], sel[2], in6[10]);
  and i107(and10[7], sel[0], sel[1], sel[2], in7[10]);

  or or10(Result[10], and10[0], and10[1], and10[2], and10[3], and10[4], and10[5], and10[6], and10[7]);

  and i110(and11[0], sel_not[0], sel_not[1], sel_not[2], in0[11]);
  and i111(and11[1], sel[0], sel_not[1], sel_not[2], in1[11]);
  and i112(and11[2], sel_not[0], sel[1], sel_not[2], in2[11]);
  and i113(and11[3], sel[0], sel[1], sel_not[2], in3[11]);
  and i114(and11[4], sel_not[0], sel_not[1], sel[2], in4[11]);
  and i115(and11[5], sel[0], sel_not[1], sel[2], in5[11]);
  and i116(and11[6], sel_not[0], sel[1], sel[2], in6[11]);
  and i117(and11[7], sel[0], sel[1], sel[2], in7[11]);

  or or11(Result[11], and11[0], and11[1], and11[2], and11[3], and11[4], and11[5], and11[6], and11[7]);

  and i120(and12[0], sel_not[0], sel_not[1], sel_not[2], in0[12]);
  and i121(and12[1], sel[0], sel_not[1], sel_not[2], in1[12]);
  and i122(and12[2], sel_not[0], sel[1], sel_not[2], in2[12]);
  and i123(and12[3], sel[0], sel[1], sel_not[2], in3[12]);
  and i124(and12[4], sel_not[0], sel_not[1], sel[2], in4[12]);
  and i125(and12[5], sel[0], sel_not[1], sel[2], in5[12]);
  and i126(and12[6], sel_not[0], sel[1], sel[2], in6[12]);
  and i127(and12[7], sel[0], sel[1], sel[2], in7[12]);

  or or12(Result[12], and12[0], and12[1], and12[2], and12[3], and12[4], and12[5], and12[6], and12[7]);

  and i130(and13[0], sel_not[0], sel_not[1], sel_not[2], in0[13]);
  and i131(and13[1], sel[0], sel_not[1], sel_not[2], in1[13]);
  and i132(and13[2], sel_not[0], sel[1], sel_not[2], in2[13]);
  and i133(and13[3], sel[0], sel[1], sel_not[2], in3[13]);
  and i134(and13[4], sel_not[0], sel_not[1], sel[2], in4[13]);
  and i135(and13[5], sel[0], sel_not[1], sel[2], in5[13]);
  and i136(and13[6], sel_not[0], sel[1], sel[2], in6[13]);
  and i137(and13[7], sel[0], sel[1], sel[2], in7[13]);

  or or13(Result[13], and13[0], and13[1], and13[2], and13[3], and13[4], and13[5], and13[6], and13[7]);

  and i140(and14[0], sel_not[0], sel_not[1], sel_not[2], in0[14]);
  and i141(and14[1], sel[0], sel_not[1], sel_not[2], in1[14]);
  and i142(and14[2], sel_not[0], sel[1], sel_not[2], in2[14]);
  and i143(and14[3], sel[0], sel[1], sel_not[2], in3[14]);
  and i144(and14[4], sel_not[0], sel_not[1], sel[2], in4[14]);
  and i145(and14[5], sel[0], sel_not[1], sel[2], in5[14]);
  and i146(and14[6], sel_not[0], sel[1], sel[2], in6[14]);
  and i147(and14[7], sel[0], sel[1], sel[2], in7[14]);

  or or14(Result[14], and14[0], and14[1], and14[2], and14[3], and14[4], and14[5], and14[6], and14[7]);

  and i150(and15[0], sel_not[0], sel_not[1], sel_not[2], in0[15]);
  and i151(and15[1], sel[0], sel_not[1], sel_not[2], in1[15]);
  and i152(and15[2], sel_not[0], sel[1], sel_not[2], in2[15]);
  and i153(and15[3], sel[0], sel[1], sel_not[2], in3[15]);
  and i154(and15[4], sel_not[0], sel_not[1], sel[2], in4[15]);
  and i155(and15[5], sel[0], sel_not[1], sel[2], in5[15]);
  and i156(and15[6], sel_not[0], sel[1], sel[2], in6[15]);
  and i157(and15[7], sel[0], sel[1], sel[2], in7[15]);

  or or15(Result[15], and15[0], and15[1], and15[2], and15[3], and15[4], and15[5], and15[6], and15[7]);

  and i160(and16[0], sel_not[0], sel_not[1], sel_not[2], in0[16]);
  and i161(and16[1], sel[0], sel_not[1], sel_not[2], in1[16]);
  and i162(and16[2], sel_not[0], sel[1], sel_not[2], in2[16]);
  and i163(and16[3], sel[0], sel[1], sel_not[2], in3[16]);
  and i164(and16[4], sel_not[0], sel_not[1], sel[2], in4[16]);
  and i165(and16[5], sel[0], sel_not[1], sel[2], in5[16]);
  and i166(and16[6], sel_not[0], sel[1], sel[2], in6[16]);
  and i167(and16[7], sel[0], sel[1], sel[2], in7[16]);

  or or16(Result[16], and16[0], and16[1], and16[2], and16[3], and16[4], and16[5], and16[6], and16[7]);

  and i170(and17[0], sel_not[0], sel_not[1], sel_not[2], in0[17]);
  and i171(and17[1], sel[0], sel_not[1], sel_not[2], in1[17]);
  and i172(and17[2], sel_not[0], sel[1], sel_not[2], in2[17]);
  and i173(and17[3], sel[0], sel[1], sel_not[2], in3[17]);
  and i174(and17[4], sel_not[0], sel_not[1], sel[2], in4[17]);
  and i175(and17[5], sel[0], sel_not[1], sel[2], in5[17]);
  and i176(and17[6], sel_not[0], sel[1], sel[2], in6[17]);
  and i177(and17[7], sel[0], sel[1], sel[2], in7[17]);

  or or17(Result[17], and17[0], and17[1], and17[2], and17[3], and17[4], and17[5], and17[6], and17[7]);

  and i180(and18[0], sel_not[0], sel_not[1], sel_not[2], in0[18]);
  and i181(and18[1], sel[0], sel_not[1], sel_not[2], in1[18]);
  and i182(and18[2], sel_not[0], sel[1], sel_not[2], in2[18]);
  and i183(and18[3], sel[0], sel[1], sel_not[2], in3[18]);
  and i184(and18[4], sel_not[0], sel_not[1], sel[2], in4[18]);
  and i185(and18[5], sel[0], sel_not[1], sel[2], in5[18]);
  and i186(and18[6], sel_not[0], sel[1], sel[2], in6[18]);
  and i187(and18[7], sel[0], sel[1], sel[2], in7[18]);

  or or18(Result[18], and18[0], and18[1], and18[2], and18[3], and18[4], and18[5], and18[6], and18[7]);

  and i190(and19[0], sel_not[0], sel_not[1], sel_not[2], in0[19]);
  and i191(and19[1], sel[0], sel_not[1], sel_not[2], in1[19]);
  and i192(and19[2], sel_not[0], sel[1], sel_not[2], in2[19]);
  and i193(and19[3], sel[0], sel[1], sel_not[2], in3[19]);
  and i194(and19[4], sel_not[0], sel_not[1], sel[2], in4[19]);
  and i195(and19[5], sel[0], sel_not[1], sel[2], in5[19]);
  and i196(and19[6], sel_not[0], sel[1], sel[2], in6[19]);
  and i197(and19[7], sel[0], sel[1], sel[2], in7[19]);

  or or19(Result[19], and19[0], and19[1], and19[2], and19[3], and19[4], and19[5], and19[6], and19[7]);

  and i200(and20[0], sel_not[0], sel_not[1], sel_not[2], in0[20]);
  and i201(and20[1], sel[0], sel_not[1], sel_not[2], in1[20]);
  and i202(and20[2], sel_not[0], sel[1], sel_not[2], in2[20]);
  and i203(and20[3], sel[0], sel[1], sel_not[2], in3[20]);
  and i204(and20[4], sel_not[0], sel_not[1], sel[2], in4[20]);
  and i205(and20[5], sel[0], sel_not[1], sel[2], in5[20]);
  and i206(and20[6], sel_not[0], sel[1], sel[2], in6[20]);
  and i207(and20[7], sel[0], sel[1], sel[2], in7[20]);

  or or20(Result[20], and20[0], and20[1], and20[2], and20[3], and20[4], and20[5], and20[6], and20[7]);

  and i210(and21[0], sel_not[0], sel_not[1], sel_not[2], in0[21]);
  and i211(and21[1], sel[0], sel_not[1], sel_not[2], in1[21]);
  and i212(and21[2], sel_not[0], sel[1], sel_not[2], in2[21]);
  and i213(and21[3], sel[0], sel[1], sel_not[2], in3[21]);
  and i214(and21[4], sel_not[0], sel_not[1], sel[2], in4[21]);
  and i215(and21[5], sel[0], sel_not[1], sel[2], in5[21]);
  and i216(and21[6], sel_not[0], sel[1], sel[2], in6[21]);
  and i217(and21[7], sel[0], sel[1], sel[2], in7[21]);

  or or21(Result[21], and21[0], and21[1], and21[2], and21[3], and21[4], and21[5], and21[6], and21[7]);

  and i220(and22[0], sel_not[0], sel_not[1], sel_not[2], in0[22]);
  and i221(and22[1], sel[0], sel_not[1], sel_not[2], in1[22]);
  and i222(and22[2], sel_not[0], sel[1], sel_not[2], in2[22]);
  and i223(and22[3], sel[0], sel[1], sel_not[2], in3[22]);
  and i224(and22[4], sel_not[0], sel_not[1], sel[2], in4[22]);
  and i225(and22[5], sel[0], sel_not[1], sel[2], in5[22]);
  and i226(and22[6], sel_not[0], sel[1], sel[2], in6[22]);
  and i227(and22[7], sel[0], sel[1], sel[2], in7[22]);

  or or22(Result[22], and22[0], and22[1], and22[2], and22[3], and22[4], and22[5], and22[6], and22[7]);

  and i230(and23[0], sel_not[0], sel_not[1], sel_not[2], in0[23]);
  and i231(and23[1], sel[0], sel_not[1], sel_not[2], in1[23]);
  and i232(and23[2], sel_not[0], sel[1], sel_not[2], in2[23]);
  and i233(and23[3], sel[0], sel[1], sel_not[2], in3[23]);
  and i234(and23[4], sel_not[0], sel_not[1], sel[2], in4[23]);
  and i235(and23[5], sel[0], sel_not[1], sel[2], in5[23]);
  and i236(and23[6], sel_not[0], sel[1], sel[2], in6[23]);
  and i237(and23[7], sel[0], sel[1], sel[2], in7[23]);

  or or23(Result[23], and23[0], and23[1], and23[2], and23[3], and23[4], and23[5], and23[6], and23[7]);

  and i240(and24[0], sel_not[0], sel_not[1], sel_not[2], in0[24]);
  and i241(and24[1], sel[0], sel_not[1], sel_not[2], in1[24]);
  and i242(and24[2], sel_not[0], sel[1], sel_not[2], in2[24]);
  and i243(and24[3], sel[0], sel[1], sel_not[2], in3[24]);
  and i244(and24[4], sel_not[0], sel_not[1], sel[2], in4[24]);
  and i245(and24[5], sel[0], sel_not[1], sel[2], in5[24]);
  and i246(and24[6], sel_not[0], sel[1], sel[2], in6[24]);
  and i247(and24[7], sel[0], sel[1], sel[2], in7[24]);

  or or24(Result[24], and24[0], and24[1], and24[2], and24[3], and24[4], and24[5], and24[6], and24[7]);

  and i250(and25[0], sel_not[0], sel_not[1], sel_not[2], in0[25]);
  and i251(and25[1], sel[0], sel_not[1], sel_not[2], in1[25]);
  and i252(and25[2], sel_not[0], sel[1], sel_not[2], in2[25]);
  and i253(and25[3], sel[0], sel[1], sel_not[2], in3[25]);
  and i254(and25[4], sel_not[0], sel_not[1], sel[2], in4[25]);
  and i255(and25[5], sel[0], sel_not[1], sel[2], in5[25]);
  and i256(and25[6], sel_not[0], sel[1], sel[2], in6[25]);
  and i257(and25[7], sel[0], sel[1], sel[2], in7[25]);

  or or25(Result[25], and25[0], and25[1], and25[2], and25[3], and25[4], and25[5], and25[6], and25[7]);

  and i260(and26[0], sel_not[0], sel_not[1], sel_not[2], in0[26]);
  and i261(and26[1], sel[0], sel_not[1], sel_not[2], in1[26]);
  and i262(and26[2], sel_not[0], sel[1], sel_not[2], in2[26]);
  and i263(and26[3], sel[0], sel[1], sel_not[2], in3[26]);
  and i264(and26[4], sel_not[0], sel_not[1], sel[2], in4[26]);
  and i265(and26[5], sel[0], sel_not[1], sel[2], in5[26]);
  and i266(and26[6], sel_not[0], sel[1], sel[2], in6[26]);
  and i267(and26[7], sel[0], sel[1], sel[2], in7[26]);

  or or26(Result[26], and26[0], and26[1], and26[2], and26[3], and26[4], and26[5], and26[6], and26[7]);

  and i270(and27[0], sel_not[0], sel_not[1], sel_not[2], in0[27]);
  and i271(and27[1], sel[0], sel_not[1], sel_not[2], in1[27]);
  and i272(and27[2], sel_not[0], sel[1], sel_not[2], in2[27]);
  and i273(and27[3], sel[0], sel[1], sel_not[2], in3[27]);
  and i274(and27[4], sel_not[0], sel_not[1], sel[2], in4[27]);
  and i275(and27[5], sel[0], sel_not[1], sel[2], in5[27]);
  and i276(and27[6], sel_not[0], sel[1], sel[2], in6[27]);
  and i277(and27[7], sel[0], sel[1], sel[2], in7[27]);

  or or27(Result[27], and27[0], and27[1], and27[2], and27[3], and27[4], and27[5], and27[6], and27[7]);

  and i280(and28[0], sel_not[0], sel_not[1], sel_not[2], in0[28]);
  and i281(and28[1], sel[0], sel_not[1], sel_not[2], in1[28]);
  and i282(and28[2], sel_not[0], sel[1], sel_not[2], in2[28]);
  and i283(and28[3], sel[0], sel[1], sel_not[2], in3[28]);
  and i284(and28[4], sel_not[0], sel_not[1], sel[2], in4[28]);
  and i285(and28[5], sel[0], sel_not[1], sel[2], in5[28]);
  and i286(and28[6], sel_not[0], sel[1], sel[2], in6[28]);
  and i287(and28[7], sel[0], sel[1], sel[2], in7[28]);

  or or28(Result[28], and28[0], and28[1], and28[2], and28[3], and28[4], and28[5], and28[6], and28[7]);

  and i290(and29[0], sel_not[0], sel_not[1], sel_not[2], in0[29]);
  and i291(and29[1], sel[0], sel_not[1], sel_not[2], in1[29]);
  and i292(and29[2], sel_not[0], sel[1], sel_not[2], in2[29]);
  and i293(and29[3], sel[0], sel[1], sel_not[2], in3[29]);
  and i294(and29[4], sel_not[0], sel_not[1], sel[2], in4[29]);
  and i295(and29[5], sel[0], sel_not[1], sel[2], in5[29]);
  and i296(and29[6], sel_not[0], sel[1], sel[2], in6[29]);
  and i297(and29[7], sel[0], sel[1], sel[2], in7[29]);

  or or29(Result[29], and29[0], and29[1], and29[2], and29[3], and29[4], and29[5], and29[6], and29[7]);

  and i300(and30[0], sel_not[0], sel_not[1], sel_not[2], in0[30]);
  and i301(and30[1], sel[0], sel_not[1], sel_not[2], in1[30]);
  and i302(and30[2], sel_not[0], sel[1], sel_not[2], in2[30]);
  and i303(and30[3], sel[0], sel[1], sel_not[2], in3[30]);
  and i304(and30[4], sel_not[0], sel_not[1], sel[2], in4[30]);
  and i305(and30[5], sel[0], sel_not[1], sel[2], in5[30]);
  and i306(and30[6], sel_not[0], sel[1], sel[2], in6[30]);
  and i307(and30[7], sel[0], sel[1], sel[2], in7[30]);

  or or30(Result[30], and30[0], and30[1], and30[2], and30[3], and30[4], and30[5], and30[6], and30[7]);

  and i310(and31[0], sel_not[0], sel_not[1], sel_not[2], in0[31]);
  and i311(and31[1], sel[0], sel_not[1], sel_not[2], in1[31]);
  and i312(and31[2], sel_not[0], sel[1], sel_not[2], in2[31]);
  and i313(and31[3], sel[0], sel[1], sel_not[2], in3[31]);
  and i314(and31[4], sel_not[0], sel_not[1], sel[2], in4[31]);
  and i315(and31[5], sel[0], sel_not[1], sel[2], in5[31]);
  and i316(and31[6], sel_not[0], sel[1], sel[2], in6[31]);
  and i317(and31[7], sel[0], sel[1], sel[2], in7[31]);

  or or31(Result[31], and31[0], and30[1], and31[2], and31[3], and31[4], and31[5], and31[6], and31[7]);

endmodule
