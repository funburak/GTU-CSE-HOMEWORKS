module and_32_bit(
	output [31:0] Result, 
	input [31:0] A,
	input [31:0] B
);

    and(Result[0], A[0], B[0]);
    and(Result[1], A[1], B[1]);
    and(Result[2], A[2], B[2]);
    and(Result[3], A[3], B[3]);
    and(Result[4], A[4], B[4]);
    and(Result[5], A[5], B[5]);
    and(Result[6], A[6], B[6]);
    and(Result[7], A[7], B[7]);
    and(Result[8], A[8], B[8]);
    and(Result[9], A[9], B[9]);
    and(Result[10], A[10], B[10]);
    and(Result[11], A[11], B[11]);
    and(Result[12], A[12], B[12]);
    and(Result[13], A[13], B[13]);
    and(Result[14], A[14], B[14]);
    and(Result[15], A[15], B[15]);
    and(Result[16], A[16], B[16]);
    and(Result[17], A[17], B[17]);
    and(Result[18], A[18], B[18]);
    and(Result[19], A[19], B[19]);
    and(Result[20], A[20], B[20]);
    and(Result[21], A[21], B[21]);
    and(Result[22], A[22], B[22]);
    and(Result[23], A[23], B[23]);
    and(Result[24], A[24], B[24]);
    and(Result[25], A[25], B[25]);
    and(Result[26], A[26], B[26]);
    and(Result[27], A[27], B[27]);
    and(Result[28], A[28], B[28]);
    and(Result[29], A[29], B[29]);
    and(Result[30], A[30], B[30]);
    and(Result[31], A[31], B[31]);

endmodule

