module not_32_bit(
	output [31:0] Result, 
	input [31:0] A
);

    not(Result[0], A[0]);
    not(Result[1], A[1]);
    not(Result[2], A[2]);
    not(Result[3], A[3]);
    not(Result[4], A[4]);
    not(Result[5], A[5]);
    not(Result[6], A[6]);
    not(Result[7], A[7]);
    not(Result[8], A[8]);
    not(Result[9], A[9]);
    not(Result[10], A[10]);
    not(Result[11], A[11]);
    not(Result[12], A[12]);
    not(Result[13], A[13]);
    not(Result[14], A[14]);
    not(Result[15], A[15]);
    not(Result[16], A[16]);
    not(Result[17], A[17]);
    not(Result[18], A[18]);
    not(Result[19], A[19]);
    not(Result[20], A[20]);
    not(Result[21], A[21]);
    not(Result[22], A[22]);
    not(Result[23], A[23]);
    not(Result[24], A[24]);
    not(Result[25], A[25]);
    not(Result[26], A[26]);
    not(Result[27], A[27]);
    not(Result[28], A[28]);
    not(Result[29], A[29]);
    not(Result[30], A[30]);
    not(Result[31], A[31]);


endmodule
