module or_32_bit(
	output [31:0] Result, 
	input [31:0] A, 
	input [31:0] B
);

    or(Result[0], A[0], B[0]);
    or(Result[1], A[1], B[1]);
    or(Result[2], A[2], B[2]);
    or(Result[3], A[3], B[3]);
    or(Result[4], A[4], B[4]);
    or(Result[5], A[5], B[5]);
    or(Result[6], A[6], B[6]);
    or(Result[7], A[7], B[7]);
    or(Result[8], A[8], B[8]);
    or(Result[9], A[9], B[9]);
    or(Result[10], A[10], B[10]);
    or(Result[11], A[11], B[11]);
    or(Result[12], A[12], B[12]);
    or(Result[13], A[13], B[13]);
    or(Result[14], A[14], B[14]);
    or(Result[15], A[15], B[15]);
    or(Result[16], A[16], B[16]);
    or(Result[17], A[17], B[17]);
    or(Result[18], A[18], B[18]);
    or(Result[19], A[19], B[19]);
    or(Result[20], A[20], B[20]);
    or(Result[21], A[21], B[21]);
    or(Result[22], A[22], B[22]);
    or(Result[23], A[23], B[23]);
    or(Result[24], A[24], B[24]);
    or(Result[25], A[25], B[25]);
    or(Result[26], A[26], B[26]);
    or(Result[27], A[27], B[27]);
    or(Result[28], A[28], B[28]);
    or(Result[29], A[29], B[29]);
    or(Result[30], A[30], B[30]);
    or(Result[31], A[31], B[31]);


endmodule
