module not_32_bit(
	input [31:0] A,
	output [31:0] Result
);

	not i0(Result[0], A[0]);
	not i1(Result[1], A[1]);
	not i2(Result[2], A[2]);
	not i3(Result[3], A[3]);
	not i4(Result[4], A[4]);
	not i5(Result[5], A[5]);
	not i6(Result[6], A[6]);
	not i7(Result[7], A[7]);
	not i8(Result[8], A[8]);
	not i9(Result[9], A[9]);
	not i10(Result[10], A[10]);
	not i11(Result[11], A[11]);
	not i12(Result[12], A[12]);
	not i13(Result[13], A[13]);
	not i14(Result[14], A[14]);
	not i15(Result[15], A[15]);
	not i16(Result[16], A[16]);
	not i17(Result[17], A[17]);
	not i18(Result[18], A[18]);
	not i19(Result[19], A[19]);
	not i20(Result[20], A[20]);
	not i21(Result[21], A[21]);
	not i22(Result[22], A[22]);
	not i23(Result[23], A[23]);
	not i24(Result[24], A[24]);
	not i25(Result[25], A[25]);
	not i26(Result[26], A[26]);
	not i27(Result[27], A[27]);
	not i28(Result[28], A[28]);
	not i29(Result[29], A[29]);
	not i30(Result[30], A[30]);
	not i31(Result[31], A[31]);



endmodule

